`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/08 17:07:05
// Design Name: 
// Module Name: tb_FA_4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_FA_4();


reg a0, a1, a2, a3, b0, b1, b2, b3, cin;
wire s0, s1, s2, s3, cout;

FA_4 dut(
    .a0(a0),
    .a1(a1),
    .a2(a2),
    .a3(a3),
    .b0(b0),
    .b1(b1),
    .b2(b2),
    .b3(b3),
    .cin(cin),
    .s0(s0),
    .s1(s1),
    .s2(s2),
    .s3(s3),
    .cout(cout)
);

initial begin 
    
    #0;
    a3 = 1'b0; a2 = 1'b0; a1 = 1'b0; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    cin = 1'b0;
    #1;//delay 값 유지
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b0; a1 = 1'b0; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b0; a1 = 1'b1; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b0; a1 = 1'b1; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b0; a0 = 1'b0;   
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b0; a0 = 1'b1;  
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b1; a0 = 1'b0;  
     b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b0; a2 = 1'b1; a1 = 1'b1; a0 = 1'b1;  
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b0; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b0; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b1; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b0; a1 = 1'b1; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b1; a1 = 1'b0; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b1; a1 = 1'b1; a0 = 1'b0;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    a3 = 1'b1; a2 = 1'b1; a1 = 1'b1; a0 = 1'b1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b0; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b0; b1 = 1'b1; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b0; b0 = 1'b1;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b0;
    #1;
    b3 = 1'b1; b2 = 1'b1; b1 = 1'b1; b0 = 1'b1;
    #1;

    $finish;



end


endmodule
