`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/15 09:37:25
// Design Name: 
// Module Name: tb_block_nonblock
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_block_nonblock();

    reg clk, a,b;
    
    initial begin
    a=0;
    b=1;
    clk=0;    
    end

    always
        clk =#5 ~clk;

    always @(posedge clk) begin
        a<=b;
        b<=a;
    end

endmodule


//////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////////////////////////////////////////////