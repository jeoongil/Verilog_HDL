`timescale 1ns / 1ps

module tb_uatr_cntl();


endmodule
