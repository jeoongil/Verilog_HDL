`timescale 1ns / 1ps

module text_practice(


    );
endmodule
